typedef struct packed {
    
} struct_floating_alu;