typedef struct packed {
    
} struct_threading_reg;