//Defining opcode and functs

//Opcode
`define Rtype 3'b000
`define Itype 3'b001
`define Mtype 3'b100
`define Ctype 3'b111
`define Ptype 3'b010
`define Xtype 3'b101

//ALUOps
`define ALU_ADD 4'b0000
`define ALU_SUB 4'b0001
`define ALU_MUL 4'b0010
`define ALU_MAC 4'b0011
`define ALU_DIV 4'b0100
`define ALU_REM 4'b0101
`define ALU_SLL 4'b0110
`define ALU_SRL 4'b0111
`define ALU_SQRT 4'b1000
`define ALU_SLT 4'b1001
`define ALU_SEQ 4'b1010
`define ALU_MAX 4'b1011
`define ALU_MIN 4'b1100
`define ALU_ABS 4'b1101
`define ALU_NOP 4'b1111

